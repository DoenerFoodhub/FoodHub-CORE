module domain

pub struct Addon {
	pub:
		id int

	pub mut:
		name string
		price f32
}