module domain

pub struct Ingredient {
	pub:
		id int

	pub mut:
		name string
		is_done bool
}