module domain

pub struct Restaurant {
	pub:
		id int

	pub mut:
		name string
		address string
		phone_number string
}